type image_matrix is array (0 to 119, 0 to 159) of std_logic_vector(11 downto 0);
constant image_data : image_matrix := (
    (