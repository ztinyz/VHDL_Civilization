type image_matrix is array (0 to 119, 0 to 159) of std_logic_vector(11 downto 0);
constant image_data : image_matrix := (
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"999", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"798", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"998", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"AA9", X"9A8", X"AA9", X"9A8", X"AA8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA9", X"9A8", X"9A8", X"AA8", X"9A8", X"AA9", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"AA9", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"8A9", X"9A9", X"9A9", X"9A9", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"AA9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA8", X"9A8", X"AA8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA9", X"AA8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA9", X"9A8", X"AA9", X"9A8", X"9A8", X"AA9", X"AA8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"898", X"898", X"898", X"898", X"898", X"AA8", X"9A8", X"AA8", X"AA9", X"AA8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"AA8", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898"),
    (X"898", X"898", X"898", X"8A9", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"AA8", X"AA9", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"AA8", X"9A8", X"AA9", X"9A8", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"998", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA9", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"8A9", X"898", X"9A9", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"8A9", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"899", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"9A9", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"9A9", X"898", X"8A8", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA8", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"AA8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"998", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A8", X"AA8", X"AA8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"8A9", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A8", X"9A8", X"AA8", X"AA8", X"9A8", X"9A8", X"AA9", X"9A8", X"AA8", X"9A8", X"9A8", X"AA8", X"9A8", X"9A8", X"9A8", X"AA8", X"9A8", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"BA8", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB9", X"AA8", X"AA8", X"BA8", X"BA8", X"898", X"898", X"898", X"998", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"8A8", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A8", X"8A9", X"8A8", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"9A8", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"8A8", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"8A9", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A9", X"898", X"898", X"898", X"9A9", X"9A9", X"898", X"8A8", X"898", X"898", X"9A9", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"8A9", X"BA8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"8A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"898"),
    (X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"AA8", X"BB8", X"9A9", X"898", X"898", X"898", X"8A9", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"999", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A8", X"898", X"998", X"898", X"898", X"898", X"898", X"9A8", X"898", X"8A8", X"898", X"9A9", X"8A8", X"898", X"898", X"9A9", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"9A8", X"8A8", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"8A8", X"898", X"898", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"BB8", X"BA8", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AB8", X"BB8", X"BA8", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A9", X"898", X"9A9", X"898", X"898", X"8A8", X"899", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"8A8", X"898", X"898", X"898", X"898", X"998", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"9A9", X"898", X"8A8", X"898", X"8A8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898"),
    (X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"998", X"898", X"898", X"898", X"898", X"9A8", X"9A9", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A8", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"9A9", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"8A8", X"898", X"9A9", X"898", X"898", X"898", X"898", X"899", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB9", X"BB8", X"BB8", X"AA8", X"BB8", X"BB8", X"BA8", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A8", X"9A9", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"898", X"8A8", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"898", X"BA8", X"BA8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"898", X"898", X"898", X"8A8", X"898", X"9A8", X"898", X"898", X"898", X"898", X"8A8", X"9A8"),
    (X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"9A8", X"898", X"898", X"8A8", X"898", X"8A8", X"9A9", X"898", X"898", X"898", X"9A9", X"898", X"898", X"9A9", X"898", X"9A8", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"AA8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"BA8", X"BB9", X"9A8", X"9A8", X"9A9", X"8A8", X"898", X"898", X"8A8", X"898", X"9A8", X"898", X"898", X"898", X"8A8", X"9A9", X"898", X"898", X"9A8", X"898", X"898", X"898", X"8A9", X"8A8", X"898", X"8A8", X"9A9", X"9A9", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"8A8", X"8A8", X"998", X"9A8", X"898", X"BA8", X"BB8", X"BB8", X"BB8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB9", X"BB9", X"898", X"898", X"998", X"898", X"9A8", X"898", X"998", X"898", X"898", X"9A9", X"9A9", X"9A9", X"898", X"9A9", X"8A8", X"898", X"898", X"898", X"898", X"8A8", X"9A8", X"898", X"9A8", X"898", X"898", X"898", X"8A8", X"9A8", X"898", X"9A8", X"9A9", X"9A8", X"898", X"9A8", X"898", X"898", X"898", X"8A9", X"898", X"9A8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"9A8", X"998", X"8A8", X"998", X"898", X"898", X"898", X"898", X"8A8", X"9A8", X"898", X"898"),
    (X"898", X"898", X"898", X"898", X"9A8", X"898", X"8A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"998", X"9A8", X"9A8", X"8A9", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"898", X"898", X"898", X"898", X"9A8", X"8A8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"8A8", X"898", X"898", X"8A8", X"898", X"9A8", X"898", X"9A9", X"9A8", X"898", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"BB8", X"BB8", X"AA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BB9", X"BA8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"898", X"8A8", X"898", X"9A8", X"9A8", X"898", X"9A8", X"8A8", X"898", X"898", X"9A8", X"898", X"9A8", X"898", X"9A9", X"8A8", X"898", X"998", X"898", X"899", X"BA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"898"),
    (X"898", X"898", X"9A9", X"9A8", X"9A8", X"8A8", X"8A8", X"898", X"898", X"9A8", X"898", X"898", X"998", X"8A8", X"9A8", X"898", X"8A8", X"9A9", X"898", X"898", X"898", X"9A8", X"9A9", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"8A8", X"898", X"898", X"898", X"898", X"8A8", X"898", X"898", X"9A8", X"898", X"9A9", X"9A8", X"898", X"9A9", X"898", X"898", X"898", X"898", X"898", X"9A8", X"8A8", X"898", X"9A8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"9A9", X"898", X"898", X"898", X"898", X"8A8", X"899", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BA8", X"898", X"9A8", X"9A8", X"898", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"9A9", X"9A9", X"898", X"9A8", X"9A8", X"898", X"898", X"898", X"9A9", X"898", X"9A9", X"898", X"898", X"899", X"BB9", X"BB8", X"BB9", X"BB8", X"BB8", X"BB9", X"CB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"CB8", X"898", X"898", X"8A8", X"898", X"8A8", X"898", X"9A8"),
    (X"898", X"9A8", X"898", X"898", X"898", X"9A8", X"898", X"9A8", X"898", X"898", X"8A8", X"9A8", X"898", X"898", X"9A8", X"898", X"898", X"898", X"898", X"9A8", X"898", X"898", X"9A9", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"9A9", X"898", X"9A8", X"9A8", X"8A8", X"9A8", X"9A9", X"898", X"9A8", X"898", X"9A8", X"898", X"998", X"9A9", X"9A8", X"898", X"9A8", X"998", X"898", X"9A8", X"898", X"898", X"898", X"898", X"898", X"899", X"8A8", X"898", X"9A8", X"898", X"9A9", X"898", X"898", X"898", X"9A8", X"998", X"898", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"9A9", X"9A9", X"9A8", X"898", X"898", X"898", X"9A8", X"9A9", X"898", X"9A8", X"898", X"898", X"998", X"8A8", X"898", X"998", X"898", X"9A8", X"898", X"9A9", X"9A9", X"898", X"8A8", X"9A8", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"8A8", X"898", X"898", X"898", X"9A9", X"898", X"9A8"),
    (X"998", X"9A9", X"898", X"8A8", X"9A8", X"998", X"9A8", X"898", X"9A9", X"898", X"898", X"9A8", X"898", X"9A8", X"998", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BA8", X"BB9", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"898", X"898", X"898", X"9A8", X"9A8", X"898", X"898", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"9A8", X"9A8", X"9A9", X"898", X"998", X"9A8", X"9A9", X"898", X"9A9", X"9A8", X"8A8", X"9A8", X"898", X"8A8", X"898", X"898", X"8A8", X"9A9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"9A9", X"9A8", X"8A8", X"9A9", X"898", X"898", X"8A8", X"998", X"998", X"9A8", X"9A9", X"898", X"898", X"9A9", X"9A9", X"9A8", X"898", X"898", X"9A8", X"9A9", X"898", X"898", X"899", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"8A8", X"898", X"898", X"9A8", X"9A8", X"9A8", X"8A8", X"898", X"9A8", X"9A9", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"AA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"8A8", X"898", X"8A8", X"9A9", X"998", X"9A8", X"898", X"899", X"BB8", X"BB8", X"AA8", X"BB9", X"BB8", X"BA8", X"BA8", X"898", X"9A9", X"8A8", X"898", X"898", X"898", X"9A8", X"9A9", X"9A8", X"898", X"9A8", X"9A8", X"9A8", X"9A9", X"898", X"8A8", X"998", X"898", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"898", X"898", X"8A8", X"9A9", X"9A8", X"9A9", X"9A8", X"898", X"998", X"898", X"9A9", X"998", X"898", X"998", X"9A8", X"998", X"8A9", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"898", X"898", X"9A8", X"898", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"898", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"898", X"8A8", X"998", X"9A9", X"9A8", X"9A9", X"898", X"8A8", X"9A8", X"9A8", X"9A8", X"9A8", X"898", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"BB8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"BA8", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"898", X"998", X"898", X"9A8", X"9A9", X"898", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"998", X"9A9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"BA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"998", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"9A8", X"9A8", X"998", X"898", X"998", X"898", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"BB9", X"BB8", X"BB8", X"BA8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"998", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"BA8", X"BB8", X"BB9", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"9A8", X"898", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"BB9", X"BB8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AB8", X"BB8", X"AA8", X"AA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"8A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"AB8", X"898", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"9A8", X"9A9", X"9A9", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BA8", X"BB8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"BA8", X"AA8", X"AA8", X"AB8", X"AA8", X"BA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"BA7", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8", X"BB8", X"BB8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8"),
    (X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"9A8", X"9A8", X"9A9", X"9A8", X"898", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9"),
    (X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"BA8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"998", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9", X"AB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"333", X"433", X"333", X"332", X"332", X"432", X"543", X"543", X"543", X"543", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"998", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"BB8", X"CCA", X"BC9", X"443", X"433", X"433", X"433", X"443", X"543", X"443", X"443", X"543", X"543", X"AB9", X"AB9", X"AB9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"998"),
    (X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BC9", X"433", X"332", X"433", X"433", X"433", X"332", X"433", X"543", X"442", X"543", X"543", X"443", X"543", X"543", X"543", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BC9", X"CCA", X"CCA", X"333", X"433", X"433", X"443", X"332", X"433", X"432", X"654", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"AB9", X"AB9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA9", X"AA9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"333", X"432", X"443", X"332", X"332", X"433", X"433", X"332", X"332", X"433", X"332", X"433", X"332", X"443", X"543", X"543", X"543", X"543", X"443", X"543", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"998", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9"),
    (X"9A8", X"AB9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"333", X"332", X"332", X"432", X"432", X"332", X"432", X"433", X"433", X"332", X"332", X"443", X"433", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"433", X"332", X"433", X"432", X"433", X"432", X"433", X"443", X"332", X"443", X"332", X"332", X"433", X"443", X"543", X"553", X"543", X"543", X"543", X"543", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"776", X"341", X"441", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"322", X"332", X"322", X"322", X"322", X"322", X"332", X"322", X"322", X"322", X"332", X"332", X"322", X"322", X"332", X"322", X"332", X"322", X"332", X"332", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"787", X"553", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"9A7", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"322", X"332", X"322", X"332", X"322", X"322", X"322", X"332", X"332", X"322", X"332", X"322", X"332", X"332", X"322", X"332", X"332", X"322", X"322", X"332", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"452", X"553", X"452", X"452", X"452", X"452", X"452", X"552", X"563", X"452", X"452", X"452", X"552", X"452", X"452", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"322", X"322", X"332", X"553", X"654", X"664", X"553", X"543", X"654", X"653", X"553", X"654", X"764", X"654", X"653", X"553", X"654", X"654", X"553", X"553", X"553", X"654", X"553", X"553", X"654", X"653", X"553", X"654", X"553", X"553", X"553", X"553", X"654", X"553", X"553", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"332", X"322", X"332", X"332", X"322", X"332", X"322", X"322", X"332", X"332", X"332", X"432", X"433", X"543", X"443", X"443", X"443", X"443", X"432", X"543", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"BB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"BB9", X"AB8", X"BA8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"452", X"562", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"553", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"322", X"332", X"322", X"664", X"654", X"653", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"653", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"553", X"554", X"653", X"553", X"553", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"332", X"322", X"322", X"322", X"322", X"322", X"332", X"332", X"322", X"332", X"433", X"443", X"433", X"443", X"443", X"443", X"543", X"442", X"543", X"543", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"BB8", X"AB8", X"AA8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9"),
    (X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"AA9", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"775", X"342", X"343", X"442", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"563", X"452", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"AB9", X"322", X"332", X"532", X"532", X"632", X"332", X"332", X"553", X"553", X"553", X"553", X"543", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"654", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"542", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"322", X"322", X"332", X"332", X"332", X"322", X"322", X"322", X"332", X"332", X"433", X"432", X"433", X"442", X"443", X"443", X"442", X"543", X"443", X"543", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"AB9", X"9A8", X"9A8", X"9A9", X"9A8", X"AA8", X"AA8", X"AB8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"BB8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8"),
    (X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AB8", X"AA8", X"AB8", X"AA8", X"AA8", X"775", X"342", X"342", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"AB9", X"322", X"332", X"532", X"633", X"632", X"332", X"332", X"654", X"664", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"664", X"553", X"553", X"553", X"543", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"542", X"AA9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"322", X"332", X"322", X"332", X"322", X"332", X"332", X"322", X"322", X"322", X"432", X"433", X"432", X"432", X"443", X"543", X"543", X"443", X"443", X"443", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"BB9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB9", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AB8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"BA8", X"9A9", X"9A9", X"342", X"342", X"443", X"342", X"443", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"342", X"342", X"452", X"452", X"452", X"452", X"452", X"452", X"442", X"552", X"AA9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"332", X"332", X"222", X"532", X"532", X"632", X"532", X"533", X"532", X"532", X"322", X"322", X"333", X"653", X"553", X"653", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"543", X"654", X"553", X"543", X"654", X"553", X"543", X"553", X"653", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"654", X"553", X"553", X"553", X"654", X"553", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"332", X"322", X"322", X"332", X"332", X"332", X"322", X"322", X"322", X"322", X"433", X"443", X"433", X"443", X"443", X"543", X"443", X"443", X"443", X"442", X"9A8", X"9A8", X"9A9", X"AB9", X"9A8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8"),
    (X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"BB8", X"9A8", X"9A9", X"342", X"342", X"342", X"342", X"342", X"452", X"563", X"664", X"452", X"452", X"563", X"452", X"563", X"342", X"342", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"552", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"322", X"322", X"332", X"532", X"632", X"633", X"632", X"532", X"532", X"532", X"322", X"322", X"322", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"664", X"553", X"553", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"654", X"553", X"553", X"553", X"553", X"765", X"553", X"553", X"654", X"654", X"553", X"553", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"332", X"322", X"322", X"322", X"322", X"332", X"322", X"332", X"322", X"332", X"332", X"433", X"443", X"432", X"443", X"443", X"443", X"443", X"543", X"543", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AB8", X"AA8", X"AA8", X"AA8", X"AA8", X"BA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB8", X"BB8"),
    (X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"AA8", X"AB8", X"AB8", X"AA8", X"AA8", X"BB9", X"CCA", X"342", X"343", X"554", X"342", X"342", X"342", X"342", X"342", X"342", X"443", X"452", X"452", X"553", X"452", X"452", X"452", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"442", X"563", X"9A9", X"9A9", X"9A8", X"9A8", X"898", X"333", X"332", X"643", X"633", X"532", X"532", X"532", X"532", X"532", X"633", X"632", X"532", X"532", X"532", X"532", X"322", X"322", X"654", X"553", X"654", X"553", X"553", X"553", X"553", X"654", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"543", X"553", X"553", X"553", X"553", X"553", X"553", X"543", X"553", X"654", X"553", X"553", X"553", X"432", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"322", X"322", X"322", X"332", X"332", X"332", X"322", X"322", X"322", X"332", X"432", X"332", X"433", X"443", X"443", X"443", X"543", X"443", X"443", X"443", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8"),
    (X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"AA8", X"BB9", X"AA8", X"AA8", X"AA8", X"BB9", X"AB9", X"AA8", X"AA8", X"CCA", X"342", X"342", X"342", X"453", X"443", X"332", X"342", X"342", X"342", X"343", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"9A9", X"9A8", X"BCA", X"BCA", X"9A8", X"544", X"322", X"532", X"633", X"532", X"532", X"632", X"532", X"632", X"532", X"643", X"532", X"532", X"532", X"643", X"322", X"322", X"553", X"553", X"553", X"553", X"553", X"553", X"654", X"553", X"653", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"554", X"653", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"543", X"442", X"ABA", X"AB9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"543", X"432", X"333", X"443", X"543", X"443", X"543", X"443", X"443", X"543", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"AA9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"AA8", X"AB9", X"AB9", X"AB8", X"AB8", X"AA8", X"AA8", X"AA8", X"AB9", X"AB8", X"AA8", X"AA8"),
    (X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A8", X"BCB", X"453", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"453", X"452", X"452", X"563", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"9A8", X"9A9", X"332", X"332", X"222", X"632", X"532", X"633", X"532", X"532", X"532", X"532", X"433", X"332", X"433", X"332", X"332", X"532", X"532", X"532", X"532", X"532", X"322", X"322", X"433", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"443", X"543", X"543", X"443", X"543", X"543", X"443", X"553", X"553", X"443", X"543", X"543", X"543", X"553", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"322", X"332", X"322", X"322", X"322", X"322", X"332", X"332", X"322", X"332", X"432", X"433", X"433", X"443", X"443", X"443", X"432", X"443", X"443", X"543", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9"),
    (X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"AA9", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"BCA", X"342", X"343", X"453", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"452", X"553", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"563", X"563", X"553", X"452", X"452", X"563", X"9A8", X"9A8", X"332", X"332", X"332", X"532", X"532", X"532", X"532", X"533", X"532", X"532", X"322", X"433", X"322", X"322", X"322", X"532", X"532", X"532", X"532", X"532", X"322", X"332", X"333", X"543", X"553", X"553", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"443", X"543", X"442", X"443", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"543", X"443", X"543", X"443", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"332", X"322", X"322", X"332", X"322", X"332", X"433", X"322", X"332", X"322", X"433", X"432", X"433", X"543", X"543", X"443", X"543", X"443", X"543", X"543", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8", X"9A8"),
    (X"9A9", X"AA9", X"9A8", X"9A9", X"9A9", X"AB9", X"9A8", X"9A9", X"9A9", X"9A8", X"AA9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"BCA", X"342", X"342", X"332", X"342", X"342", X"342", X"342", X"342", X"443", X"342", X"342", X"443", X"452", X"452", X"452", X"342", X"342", X"443", X"342", X"453", X"452", X"452", X"452", X"452", X"562", X"AA9", X"9A9", X"221", X"332", X"322", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"332", X"332", X"322", X"322", X"332", X"532", X"632", X"532", X"532", X"532", X"322", X"322", X"332", X"543", X"543", X"543", X"543", X"553", X"543", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"443", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"443", X"543", X"543", X"543", X"543", X"9A9", X"9A8", X"AA9", X"9A9", X"9A8", X"322", X"322", X"322", X"322", X"332", X"332", X"433", X"332", X"322", X"322", X"433", X"432", X"332", X"543", X"432", X"432", X"442", X"443", X"543", X"443", X"9A8", X"9A8", X"9A9", X"9A9", X"AA9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"AA9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A8", X"AA9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A9"),
    (X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"AA9", X"AA9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"AA9", X"9A9", X"9A9", X"9A9", X"9A8", X"BCA", X"342", X"342", X"332", X"342", X"342", X"342", X"342", X"342", X"342", X"343", X"342", X"443", X"342", X"342", X"342", X"342", X"342", X"332", X"443", X"453", X"442", X"452", X"452", X"452", X"451", X"332", X"332", X"633", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"633", X"643", X"633", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"633", X"532", X"532", X"332", X"322", X"543", X"543", X"553", X"442", X"543", X"543", X"443", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"443", X"553", X"9A8", X"9A9", X"322", X"322", X"322", X"322", X"332", X"322", X"322", X"322", X"322", X"322", X"433", X"443", X"433", X"443", X"432", X"332", X"332", X"322", X"543", X"553", X"553", X"553", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"654", X"553", X"553", X"553", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A9"),
    (X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"AA9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"AA9", X"BCB", X"342", X"453", X"443", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"453", X"452", X"452", X"452", X"452", X"462", X"322", X"332", X"532", X"632", X"532", X"532", X"532", X"532", X"633", X"532", X"532", X"643", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"332", X"332", X"543", X"443", X"543", X"543", X"543", X"543", X"443", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"543", X"443", X"553", X"653", X"9A8", X"9A8", X"322", X"332", X"322", X"322", X"332", X"332", X"332", X"322", X"332", X"332", X"332", X"433", X"332", X"442", X"442", X"332", X"322", X"332", X"654", X"654", X"553", X"553", X"664", X"553", X"553", X"553", X"653", X"553", X"553", X"553", X"553", X"654", X"553", X"553", X"553", X"9A8", X"9A8", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"AA9", X"9A9", X"9A9", X"9A9", X"9A9", X"AA9", X"9A9", X"9A8"),
    (X"9A9", X"9A9", X"9A8", X"9A9", X"AA9", X"9A9", X"9A9", X"9A9", X"AA9", X"9A8", X"AA9", X"9A9", X"AA9", X"AA9", X"9A8", X"9A9", X"AA9", X"AA9", X"9A9", X"9A8", X"342", X"342", X"342", X"342", X"342", X"342", X"332", X"443", X"342", X"342", X"342", X"342", X"342", X"342", X"343", X"342", X"342", X"342", X"342", X"342", X"433", X"322", X"332", X"643", X"532", X"532", X"633", X"532", X"643", X"633", X"532", X"532", X"532", X"532", X"632", X"532", X"633", X"532", X"532", X"532", X"633", X"532", X"532", X"532", X"532", X"532", X"532", X"632", X"322", X"332", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"443", X"654", X"543", X"543", X"553", X"543", X"543", X"543", X"543", X"443", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"9A9", X"9A8", X"322", X"322", X"332", X"332", X"322", X"433", X"433", X"322", X"322", X"322", X"433", X"433", X"433", X"322", X"332", X"443", X"432", X"543", X"333", X"332", X"553", X"553", X"553", X"653", X"653", X"553", X"553", X"553", X"654", X"553", X"553", X"553", X"553", X"654", X"553", X"543", X"553", X"654", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"9A8", X"AA9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"AA9", X"9A9", X"9A8"),
    (X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"AA9", X"9A9", X"AA9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A9", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"AA9", X"9A8", X"342", X"453", X"342", X"343", X"342", X"342", X"342", X"443", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"322", X"322", X"333", X"532", X"532", X"643", X"532", X"532", X"532", X"532", X"532", X"643", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"643", X"532", X"532", X"532", X"532", X"532", X"532", X"332", X"322", X"543", X"443", X"443", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"543", X"553", X"543", X"553", X"543", X"543", X"543", X"543", X"543", X"653", X"9A8", X"9A8", X"332", X"332", X"332", X"322", X"332", X"322", X"322", X"322", X"322", X"322", X"433", X"443", X"433", X"322", X"433", X"433", X"432", X"543", X"322", X"322", X"553", X"653", X"653", X"553", X"553", X"553", X"553", X"653", X"553", X"654", X"553", X"553", X"553", X"653", X"654", X"553", X"553", X"764", X"AA9", X"9A9", X"9A8", X"9A9", X"AA9", X"9A9", X"9A8", X"9A8", X"9A8", X"AB9", X"9A9", X"9A8", X"9A9", X"9A8", X"9A9", X"9A9", X"9A9"),
    (X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"553", X"453", X"453", X"9A8", X"9A9", X"9A8", X"9A9", X"9A8", X"AA9", X"AA9", X"9A8", X"342", X"343", X"342", X"443", X"342", X"342", X"342", X"342", X"332", X"342", X"443", X"342", X"342", X"554", X"342", X"342", X"342", X"342", X"332", X"342", X"9A8", X"9A8", X"9A9", X"532", X"532", X"532", X"532", X"532", X"632", X"532", X"532", X"633", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"633", X"532", X"532", X"643", X"633", X"643", X"532", X"522", X"522", X"422", X"532", X"522", X"422", X"533", X"522", X"422", X"422", X"522", X"522", X"422", X"532", X"532", X"522", X"422", X"522", X"522", X"522", X"533", X"522", X"422", X"522", X"422", X"522", X"522", X"522", X"522", X"522", X"522", X"532", X"533", X"9A8", X"9A8", X"322", X"322", X"322", X"322", X"322", X"322", X"332", X"433", X"332", X"322", X"322", X"332", X"322", X"432", X"443", X"443", X"443", X"543", X"543", X"543", X"332", X"322", X"322", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"553", X"553", X"653", X"653", X"653", X"553", X"653", X"654", X"9A8", X"9A9", X"9A8", X"9A8", X"9A9", X"9A8", X"9A8", X"ABA", X"453", X"453", X"553", X"564", X"453", X"453", X"564"),
    (X"453", X"442", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"AA9", X"9A9", X"9A9", X"AA9", X"9A9", X"9A9", X"9A8", X"9A8", X"342", X"342", X"342", X"443", X"443", X"332", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"343", X"342", X"443", X"453", X"342", X"AA9", X"9A9", X"9B9", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"632", X"532", X"532", X"532", X"632", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"643", X"532", X"532", X"643", X"532", X"532", X"532", X"422", X"422", X"522", X"421", X"532", X"522", X"532", X"422", X"422", X"532", X"522", X"422", X"422", X"522", X"422", X"532", X"422", X"522", X"522", X"522", X"422", X"522", X"421", X"522", X"522", X"422", X"532", X"422", X"522", X"522", X"522", X"9A8", X"9A9", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"322", X"332", X"322", X"322", X"332", X"333", X"443", X"443", X"443", X"442", X"432", X"432", X"443", X"322", X"332", X"222", X"653", X"664", X"553", X"654", X"553", X"553", X"553", X"553", X"553", X"553", X"653", X"553", X"553", X"553", X"553", X"553", X"653", X"AA8", X"9A8", X"9A8", X"9A9", X"9A9", X"9A8", X"9A9", X"BBA", X"453", X"453", X"453", X"453", X"453", X"453", X"453"),
    (X"453", X"342", X"453", X"453", X"564", X"553", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"564", X"453", X"343", X"453", X"564", X"443", X"453", X"453", X"453", X"342", X"342", X"342", X"453", X"343", X"343", X"332", X"332", X"342", X"342", X"342", X"342", X"342", X"453", X"342", X"AB9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"532", X"532", X"532", X"633", X"532", X"532", X"532", X"332", X"322", X"322", X"322", X"322", X"322", X"332", X"432", X"322", X"322", X"332", X"332", X"333", X"532", X"532", X"532", X"633", X"643", X"532", X"633", X"632", X"743", X"743", X"632", X"743", X"642", X"743", X"642", X"632", X"642", X"743", X"643", X"632", X"743", X"642", X"642", X"854", X"632", X"743", X"632", X"743", X"642", X"632", X"743", X"743", X"642", X"743", X"743", X"642", X"743", X"642", X"642", X"843", X"9A8", X"9A8", X"332", X"322", X"433", X"322", X"322", X"322", X"322", X"332", X"322", X"322", X"443", X"432", X"432", X"543", X"443", X"432", X"442", X"432", X"443", X"433", X"443", X"443", X"432", X"433", X"332", X"653", X"653", X"553", X"654", X"553", X"553", X"553", X"764", X"553", X"654", X"553", X"653", X"553", X"553", X"653", X"553", X"653", X"553", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453"),
    (X"453", X"553", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"564", X"342", X"342", X"342", X"342", X"443", X"342", X"322", X"332", X"342", X"342", X"342", X"342", X"332", X"342", X"342", X"AB9", X"9A9", X"9A8", X"9A8", X"9A8", X"9A9", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"332", X"332", X"332", X"433", X"322", X"322", X"332", X"322", X"332", X"332", X"322", X"322", X"222", X"532", X"632", X"532", X"532", X"532", X"532", X"532", X"632", X"743", X"632", X"743", X"743", X"743", X"743", X"632", X"742", X"632", X"742", X"742", X"643", X"743", X"743", X"743", X"743", X"632", X"743", X"743", X"743", X"742", X"642", X"742", X"632", X"632", X"743", X"742", X"743", X"632", X"743", X"642", X"743", X"9A8", X"9A8", X"322", X"322", X"433", X"332", X"322", X"332", X"332", X"433", X"332", X"332", X"543", X"432", X"443", X"543", X"543", X"432", X"442", X"443", X"443", X"443", X"442", X"443", X"432", X"433", X"332", X"553", X"553", X"653", X"654", X"653", X"553", X"553", X"553", X"553", X"553", X"654", X"553", X"553", X"653", X"553", X"654", X"553", X"643", X"443", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453"),
    (X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"454", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"342", X"322", X"332", X"332", X"322", X"332", X"332", X"332", X"453", X"453", X"443", X"453", X"453", X"564", X"453", X"453", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"322", X"332", X"322", X"322", X"332", X"322", X"332", X"332", X"322", X"322", X"322", X"322", X"222", X"532", X"532", X"633", X"532", X"532", X"532", X"643", X"743", X"743", X"642", X"743", X"742", X"642", X"643", X"732", X"322", X"332", X"743", X"743", X"743", X"642", X"743", X"743", X"743", X"742", X"322", X"332", X"742", X"743", X"632", X"743", X"642", X"632", X"743", X"632", X"743", X"743", X"632", X"642", X"732", X"453", X"453", X"322", X"332", X"322", X"332", X"322", X"332", X"332", X"322", X"443", X"432", X"432", X"443", X"442", X"432", X"443", X"543", X"543", X"443", X"443", X"442", X"443", X"443", X"443", X"543", X"433", X"443", X"432", X"543", X"443", X"443", X"543", X"442", X"443", X"543", X"443", X"543", X"443", X"443", X"443", X"443", X"443", X"442", X"543", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"564", X"453", X"453", X"453", X"453"),
    (X"453", X"453", X"453", X"453", X"453", X"452", X"453", X"452", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"553", X"453", X"453", X"453", X"453", X"453", X"342", X"332", X"433", X"322", X"443", X"332", X"322", X"332", X"453", X"453", X"453", X"564", X"453", X"453", X"453", X"353", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"322", X"332", X"322", X"332", X"322", X"433", X"322", X"332", X"322", X"332", X"332", X"322", X"332", X"532", X"532", X"532", X"633", X"632", X"532", X"532", X"743", X"743", X"642", X"742", X"743", X"642", X"632", X"954", X"322", X"332", X"632", X"642", X"632", X"743", X"632", X"743", X"632", X"632", X"332", X"322", X"743", X"632", X"732", X"743", X"743", X"742", X"742", X"743", X"632", X"743", X"743", X"743", X"732", X"453", X"453", X"322", X"332", X"433", X"322", X"322", X"332", X"322", X"332", X"443", X"432", X"432", X"433", X"443", X"543", X"432", X"433", X"443", X"433", X"443", X"443", X"442", X"432", X"443", X"443", X"543", X"543", X"443", X"443", X"442", X"543", X"432", X"442", X"443", X"443", X"543", X"543", X"443", X"443", X"443", X"443", X"443", X"442", X"543", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453"),
    (X"453", X"453", X"453", X"343", X"443", X"342", X"342", X"343", X"342", X"342", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"443", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"443", X"453", X"453", X"322", X"332", X"332", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"353", X"532", X"532", X"532", X"632", X"532", X"532", X"532", X"322", X"322", X"322", X"332", X"433", X"332", X"322", X"332", X"322", X"322", X"322", X"332", X"333", X"532", X"532", X"532", X"532", X"532", X"532", X"532", X"743", X"742", X"642", X"642", X"642", X"742", X"632", X"843", X"322", X"322", X"742", X"642", X"632", X"742", X"742", X"632", X"743", X"632", X"322", X"322", X"743", X"642", X"742", X"642", X"732", X"743", X"743", X"743", X"643", X"642", X"642", X"743", X"742", X"453", X"453", X"322", X"332", X"332", X"332", X"332", X"322", X"332", X"322", X"443", X"543", X"432", X"432", X"543", X"332", X"332", X"332", X"332", X"333", X"443", X"443", X"543", X"443", X"443", X"443", X"543", X"553", X"653", X"653", X"654", X"553", X"543", X"443", X"543", X"332", X"322", X"543", X"653", X"653", X"654", X"543", X"543", X"654", X"653", X"442", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453"),
    (X"453", X"453", X"453", X"342", X"343", X"343", X"342", X"443", X"443", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"442", X"453", X"322", X"332", X"332", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"343", X"643", X"532", X"532", X"643", X"532", X"532", X"532", X"322", X"322", X"332", X"332", X"332", X"332", X"332", X"322", X"322", X"322", X"332", X"322", X"332", X"532", X"643", X"532", X"532", X"532", X"532", X"532", X"743", X"743", X"743", X"642", X"742", X"742", X"743", X"742", X"322", X"443", X"743", X"743", X"743", X"742", X"743", X"642", X"642", X"743", X"222", X"332", X"742", X"743", X"743", X"743", X"743", X"743", X"743", X"642", X"743", X"743", X"743", X"743", X"732", X"453", X"453", X"322", X"332", X"322", X"322", X"322", X"322", X"332", X"322", X"443", X"432", X"443", X"443", X"543", X"322", X"332", X"332", X"322", X"332", X"543", X"443", X"543", X"443", X"543", X"543", X"432", X"553", X"654", X"553", X"653", X"553", X"432", X"443", X"543", X"322", X"322", X"653", X"653", X"653", X"543", X"653", X"553", X"543", X"653", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"452", X"564", X"453", X"453"),
    (X"453", X"342", X"342", X"343", X"342", X"443", X"342", X"443", X"342", X"443", X"343", X"342", X"342", X"343", X"342", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"564", X"453", X"453", X"442", X"322", X"322", X"332", X"553", X"563", X"453", X"453", X"342", X"342", X"342", X"342", X"342", X"342", X"532", X"532", X"532", X"643", X"532", X"532", X"532", X"332", X"332", X"332", X"332", X"322", X"332", X"322", X"332", X"332", X"332", X"322", X"332", X"332", X"532", X"532", X"633", X"633", X"532", X"643", X"532", X"742", X"743", X"743", X"743", X"743", X"642", X"853", X"642", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"642", X"743", X"642", X"743", X"743", X"743", X"743", X"743", X"742", X"743", X"853", X"632", X"632", X"642", X"743", X"743", X"732", X"453", X"342", X"322", X"332", X"322", X"322", X"322", X"322", X"322", X"332", X"443", X"443", X"442", X"443", X"543", X"332", X"322", X"322", X"332", X"322", X"543", X"443", X"443", X"554", X"543", X"543", X"443", X"553", X"653", X"653", X"754", X"653", X"443", X"442", X"543", X"332", X"332", X"653", X"654", X"653", X"653", X"653", X"653", X"653", X"653", X"453", X"443", X"453", X"453", X"443", X"342", X"342", X"343", X"342", X"343", X"342", X"453"),
    (X"342", X"343", X"342", X"342", X"453", X"554", X"342", X"443", X"342", X"342", X"343", X"342", X"342", X"342", X"342", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"453", X"564", X"453", X"443", X"342", X"453", X"453", X"332", X"332", X"332", X"453", X"343", X"342", X"343", X"453", X"342", X"343", X"342", X"342", X"243", X"532", X"532", X"532", X"632", X"532", X"632", X"532", X"332", X"332", X"332", X"322", X"332", X"332", X"332", X"322", X"322", X"332", X"322", X"332", X"333", X"532", X"643", X"632", X"532", X"632", X"532", X"532", X"743", X"742", X"742", X"642", X"642", X"732", X"743", X"632", X"743", X"743", X"743", X"743", X"742", X"743", X"743", X"743", X"742", X"743", X"632", X"632", X"743", X"743", X"743", X"632", X"743", X"854", X"742", X"743", X"743", X"742", X"743", X"632", X"732", X"343", X"342", X"332", X"322", X"332", X"322", X"322", X"322", X"322", X"322", X"443", X"543", X"543", X"443", X"442", X"322", X"322", X"322", X"332", X"322", X"443", X"432", X"443", X"543", X"432", X"442", X"443", X"543", X"553", X"653", X"654", X"653", X"653", X"543", X"543", X"443", X"443", X"653", X"553", X"653", X"653", X"653", X"653", X"653", X"643", X"453", X"453", X"453", X"453", X"453", X"342", X"443", X"343", X"342", X"342", X"342", X"453"),
    (X"342", X"342", X"332", X"342", X"342", X"342", X"342", X"443", X"342", X"342", X"342", X"443", X"343", X"342", X"343", X"343", X"342", X"342", X"342", X"343", X"443", X"343", X"453", X"554", X"453", X"342", X"454", X"342", X"342", X"342", X"332", X"322", X"322", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"342", X"343", X"232", X"633", X"632", X"522", X"532", X"532", X"633", X"532", X"332", X"322", X"332", X"322", X"332", X"332", X"332", X"433", X"332", X"322", X"332", X"332", X"332", X"632", X"532", X"532", X"532", X"532", X"532", X"532", X"742", X"743", X"743", X"742", X"642", X"743", X"743", X"743", X"743", X"743", X"742", X"743", X"743", X"743", X"743", X"632", X"743", X"642", X"743", X"743", X"742", X"642", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"743", X"843", X"453", X"342", X"322", X"322", X"322", X"322", X"322", X"322", X"332", X"332", X"543", X"443", X"443", X"432", X"443", X"332", X"332", X"433", X"332", X"322", X"443", X"443", X"443", X"543", X"443", X"443", X"543", X"653", X"653", X"653", X"653", X"553", X"553", X"653", X"653", X"653", X"653", X"654", X"653", X"654", X"653", X"653", X"653", X"653", X"643", X"343", X"443", X"443", X"342", X"443", X"342", X"342", X"342", X"342", X"342", X"342", X"342"),
    (X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"552", X"552", X"552", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"552", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"563", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"663", X"662", X"562", X"673", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"552", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562"),
    (X"562", X"562", X"663", X"663", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"552", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"552", X"663", X"562", X"552", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"673", X"562", X"562", X"562", X"562", X"663", X"663", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"663", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562"),
    (X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"673", X"562", X"662", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"563", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"663", X"562", X"552", X"562", X"662", X"562", X"663", X"562", X"673", X"562", X"552", X"562", X"562", X"663", X"562", X"562", X"663", X"562", X"662", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"773", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562"),
    (X"562", X"562", X"562", X"663", X"562", X"562", X"662", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"662", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"552", X"562", X"663", X"662", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"662", X"562", X"552", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562"),
    (X"562", X"562", X"562", X"562", X"663", X"662", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"663", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"662", X"562", X"662", X"562", X"562", X"673", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"772", X"772", X"773", X"773", X"772", X"772", X"772", X"772", X"772", X"772", X"773", X"773", X"772", X"773", X"873", X"773", X"773", X"873", X"873", X"772", X"772", X"772", X"873", X"773", X"772", X"772", X"772", X"883", X"773", X"772", X"873", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"A83", X"983"),
    (X"562", X"663", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"663", X"562", X"673", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"772", X"873", X"773", X"873", X"772", X"772", X"772", X"773", X"773", X"773", X"772", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"873", X"772", X"873", X"873", X"773", X"773", X"772", X"873", X"772", X"773", X"772", X"772", X"772", X"772", X"773", X"983", X"983", X"983", X"983", X"994", X"983", X"A94"),
    (X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"552", X"552", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"552", X"452", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"441", X"452", X"452", X"563", X"563", X"452", X"452", X"563", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"562", X"552", X"552", X"673", X"883", X"773", X"773", X"772", X"772", X"773", X"772", X"873", X"773", X"772", X"772", X"772", X"772", X"772", X"772", X"772", X"773", X"772", X"772", X"772", X"773", X"772", X"873", X"773", X"772", X"983", X"983", X"A94", X"983", X"A84", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"873", X"873", X"772", X"773", X"773", X"772", X"772", X"772", X"772", X"773", X"873", X"873", X"873", X"873"),
    (X"452", X"452", X"452", X"552", X"552", X"563", X"552", X"452", X"452", X"452", X"452", X"562", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"562", X"673", X"562", X"552", X"662", X"562", X"662", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"563", X"452", X"452", X"452", X"563", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"552", X"563", X"452", X"452", X"552", X"452", X"552", X"562", X"552", X"663", X"873", X"773", X"773", X"773", X"773", X"773", X"772", X"883", X"773", X"773", X"873", X"873", X"773", X"772", X"773", X"773", X"772", X"772", X"772", X"772", X"883", X"773", X"772", X"873", X"662", X"983", X"983", X"A84", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"772", X"772", X"873", X"772", X"772", X"773", X"773", X"773", X"772", X"772", X"772", X"773"),
    (X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"662", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"662", X"662", X"673", X"662", X"662", X"562", X"662", X"773", X"772", X"772", X"873", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"984", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"873", X"773", X"773", X"873", X"883", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"983", X"983", X"A94", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983"),
    (X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"662", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"552", X"452", X"562", X"452", X"552", X"552", X"563", X"452", X"452", X"452", X"562", X"552", X"452", X"452", X"773", X"662", X"662", X"662", X"552", X"662", X"662", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"A83", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"A94", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"873", X"772", X"773", X"772", X"772", X"772", X"773", X"984", X"772", X"773", X"773", X"772", X"772", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"994", X"983", X"983", X"983", X"983"),
    (X"562", X"562", X"562", X"663", X"562", X"562", X"773", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"663", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"552", X"452", X"552", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"552", X"563", X"452", X"662", X"673", X"662", X"662", X"773", X"673", X"662", X"884", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"A94", X"772", X"772", X"773", X"772", X"773", X"873", X"773", X"773", X"773", X"773", X"772", X"873", X"772", X"773", X"773", X"772", X"772", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"772", X"772", X"773", X"883", X"773", X"772", X"773", X"772", X"773", X"873", X"772", X"773", X"873", X"773", X"773", X"772", X"772", X"773", X"884", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"662", X"562", X"562", X"562", X"662", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"672", X"562", X"562", X"562", X"452", X"452", X"552", X"552", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"453", X"442", X"453", X"452", X"453", X"452", X"452", X"342", X"452", X"662", X"662", X"652", X"662", X"662", X"663", X"662", X"662", X"A93", X"A93", X"A93", X"993", X"A94", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"873", X"773", X"773", X"772", X"773", X"773", X"873", X"773", X"A93", X"A93", X"A94", X"A94", X"A94", X"A93", X"A93", X"A93", X"983", X"A94", X"A94", X"983", X"A83", X"A94", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"A83", X"883", X"773", X"773", X"773", X"773", X"783", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"772", X"773", X"873", X"883", X"983", X"A93", X"A94", X"A94", X"A93", X"A83", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983"),
    (X"452", X"563", X"452", X"452", X"563", X"563", X"452", X"552", X"552", X"552", X"563", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"662", X"663", X"562", X"663", X"673", X"663", X"662", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"662", X"673", X"993", X"983", X"983", X"983", X"A94", X"A94", X"993", X"983", X"983", X"983", X"772", X"873", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"772", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"773", X"883", X"773", X"772", X"873", X"772", X"773", X"773", X"773", X"772", X"773", X"772", X"773", X"873", X"773", X"773", X"772", X"773", X"772", X"772", X"773", X"772", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"A83", X"772", X"772", X"772", X"772", X"773", X"873", X"772", X"772", X"773", X"772", X"873", X"772", X"772", X"773", X"773", X"773", X"773", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"562", X"662", X"562", X"562", X"562", X"662", X"673", X"662", X"562", X"662", X"662", X"562", X"663", X"663", X"662", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"330", X"341", X"341", X"341", X"341", X"341", X"441", X"441", X"441", X"452", X"662", X"662", X"983", X"994", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"762", X"772", X"772", X"772", X"772", X"772", X"883", X"772", X"772", X"883", X"773", X"772", X"773", X"A94", X"A94", X"A93", X"A94", X"993", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"772", X"762", X"772", X"772", X"772", X"772", X"772", X"762", X"772", X"772", X"773", X"883", X"773", X"773", X"773", X"773", X"773", X"883", X"772", X"773", X"772", X"773", X"A94", X"993", X"983", X"983", X"983", X"993", X"A94", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"772", X"772", X"772", X"662", X"873", X"883", X"773", X"883", X"773", X"772", X"773", X"772", X"772", X"772", X"983", X"993", X"983", X"A94", X"983", X"A94", X"A94", X"A94", X"A94", X"A94"),
    (X"562", X"562", X"562", X"673", X"562", X"562", X"662", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"552", X"452", X"452", X"452", X"552", X"552", X"452", X"563", X"452", X"562", X"452", X"452", X"552", X"552", X"452", X"452", X"563", X"552", X"552", X"452", X"452", X"452", X"452", X"984", X"983", X"983", X"A94", X"983", X"983", X"A83", X"773", X"773", X"772", X"773", X"772", X"773", X"772", X"772", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"772", X"772", X"772", X"772", X"772", X"773", X"773", X"883", X"772", X"873", X"773", X"772", X"A93", X"983", X"A94", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"A94", X"983", X"873", X"773", X"772", X"773", X"772", X"773", X"873", X"883", X"883", X"772", X"772", X"873", X"883", X"773", X"883", X"773", X"772", X"773", X"773", X"773", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"773", X"772", X"772", X"873", X"772", X"773", X"773", X"773", X"873", X"883", X"772", X"773", X"773", X"873", X"772", X"873", X"772", X"773", X"773", X"773"),
    (X"673", X"562", X"662", X"562", X"562", X"451", X"552", X"452", X"452", X"452", X"452", X"451", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"563", X"662", X"663", X"662", X"662", X"773", X"773", X"773", X"873", X"773", X"883", X"873", X"873", X"873", X"873", X"873", X"883", X"773", X"993", X"993", X"983", X"983", X"993", X"A94", X"A94", X"983", X"772", X"773", X"773", X"773", X"883", X"773", X"873", X"773", X"773", X"772", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"A83", X"993", X"983", X"983", X"983", X"773", X"772", X"873", X"772", X"773", X"772", X"773", X"773", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"A94", X"983", X"A93", X"993", X"993", X"983", X"A83", X"873", X"772", X"772", X"873", X"873", X"772", X"772", X"773", X"772", X"873", X"773", X"883", X"772", X"772", X"773", X"773", X"873", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"A94", X"983", X"A93", X"983", X"984", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"773", X"772", X"772", X"773", X"772", X"773", X"773", X"772", X"772", X"773"),
    (X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"563", X"563", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"662", X"662", X"662", X"662", X"662", X"873", X"772", X"773", X"873", X"772", X"772", X"772", X"773", X"773", X"773", X"883", X"773", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"A93", X"772", X"773", X"773", X"773", X"873", X"772", X"773", X"773", X"883", X"873", X"772", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"772", X"773", X"772", X"873", X"773", X"773", X"773", X"873", X"772", X"873", X"773", X"773", X"772", X"873", X"773", X"772", X"883", X"993", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"772", X"773", X"883", X"773", X"873", X"773", X"873", X"773", X"773", X"772", X"772", X"772", X"873", X"873", X"772", X"773", X"772", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"772", X"772", X"773", X"773", X"873", X"772", X"772", X"773", X"883", X"772", X"772"),
    (X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"873", X"883", X"873", X"873", X"883", X"873", X"873", X"873", X"A94", X"A94", X"A94", X"983", X"A93", X"A94", X"983", X"993", X"983", X"A83", X"883", X"773", X"873", X"773", X"772", X"773", X"772", X"873", X"773", X"772", X"983", X"994", X"983", X"983", X"983", X"A93", X"A94", X"983", X"A94", X"A94", X"873", X"773", X"772", X"772", X"773", X"773", X"772", X"883", X"773", X"772", X"873", X"772", X"993", X"983", X"983", X"983", X"983", X"A94", X"983", X"A94", X"A94", X"A94", X"873", X"772", X"773", X"772", X"772", X"773", X"873", X"883", X"773", X"773", X"773", X"772", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"A94", X"983", X"A83", X"A93", X"983", X"993", X"983", X"983", X"983", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"772", X"772", X"773", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"984", X"993", X"A94", X"A93", X"983", X"993", X"A94", X"883", X"772", X"773", X"883", X"773"),
    (X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"563", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"873", X"772", X"772", X"772", X"773", X"773", X"773", X"773", X"993", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"772", X"773", X"773", X"773", X"873", X"873", X"773", X"883", X"772", X"773", X"983", X"A94", X"983", X"993", X"983", X"983", X"983", X"993", X"983", X"983", X"773", X"773", X"773", X"772", X"873", X"773", X"873", X"873", X"773", X"773", X"773", X"773", X"A94", X"993", X"993", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"773", X"773", X"883", X"773", X"773", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"873", X"873", X"772", X"873", X"772", X"772", X"772", X"983", X"A94", X"983", X"A94", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"873", X"772", X"873", X"773", X"873", X"773", X"883", X"772", X"772", X"883", X"772", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"883", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"A83", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"A94", X"983", X"983", X"983", X"983", X"772", X"773", X"773", X"773", X"773"),
    (X"452", X"452", X"452", X"452", X"553", X"873", X"873", X"772", X"772", X"873", X"983", X"983", X"983", X"983", X"983", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"873", X"873", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"873", X"773", X"873", X"773", X"873", X"773", X"773", X"873", X"873", X"773", X"772", X"773", X"773", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"883", X"772", X"773", X"873", X"773", X"773", X"873", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"873", X"772", X"773", X"772", X"773", X"772", X"772", X"773", X"772", X"772", X"873", X"773", X"773", X"772", X"773", X"773", X"772", X"773", X"772", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"873", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"772", X"883", X"772", X"773", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"552", X"452", X"552", X"452", X"452", X"773", X"773", X"873", X"772", X"773", X"983", X"A94", X"A94", X"983", X"983", X"873", X"773", X"773", X"873", X"773", X"773", X"772", X"873", X"873", X"773", X"983", X"983", X"983", X"983", X"A93", X"A94", X"993", X"983", X"983", X"983", X"873", X"773", X"772", X"873", X"773", X"773", X"772", X"773", X"873", X"773", X"773", X"772", X"772", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"772", X"773", X"873", X"883", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"A83", X"873", X"772", X"873", X"773", X"883", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"772", X"773", X"873", X"773", X"772", X"772", X"773", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"993", X"983", X"983", X"983", X"983", X"993", X"A94", X"983", X"A93", X"772", X"773", X"772", X"773", X"873", X"773", X"873", X"773", X"773", X"772", X"773", X"873", X"772", X"884", X"772", X"772", X"773", X"773", X"772", X"884", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"994", X"983", X"983", X"983", X"983"),
    (X"773", X"773", X"873", X"773", X"773", X"773", X"873", X"773", X"773", X"773", X"983", X"983", X"A94", X"983", X"983", X"983", X"A94", X"A83", X"773", X"773", X"773", X"773", X"772", X"772", X"873", X"873", X"773", X"884", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"773", X"873", X"873", X"773", X"772", X"772", X"773", X"873", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"984", X"993", X"983", X"983", X"983", X"773", X"772", X"772", X"773", X"772", X"873", X"873", X"772", X"773", X"773", X"873", X"772", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"993", X"994", X"983", X"773", X"772", X"873", X"773", X"772", X"883", X"772", X"773", X"773", X"873", X"773", X"772", X"773", X"883", X"772", X"773", X"873", X"772", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"873", X"883", X"773", X"773", X"772", X"772", X"772", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"772", X"773", X"772", X"772", X"873", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983"),
    (X"773", X"873", X"773", X"772", X"773", X"772", X"883", X"873", X"883", X"873", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"773", X"773", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"994", X"983", X"983", X"983", X"993", X"983", X"773", X"873", X"772", X"773", X"772", X"773", X"873", X"772", X"883", X"772", X"772", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"873", X"772", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"873", X"773", X"993", X"983", X"A94", X"A94", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"772", X"773", X"772", X"772", X"873", X"772", X"873", X"773", X"773", X"773", X"773", X"873", X"983", X"A94", X"983", X"983", X"983", X"994", X"983", X"984", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"773", X"873", X"773", X"873", X"873", X"773", X"772", X"772", X"873", X"773", X"772", X"772", X"773", X"883", X"773", X"883", X"773", X"773", X"773", X"773", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"773", X"773", X"873", X"883", X"772", X"773", X"773", X"873", X"773", X"873", X"873", X"772", X"883", X"A94", X"983", X"983", X"983", X"983", X"873", X"873", X"773", X"773", X"773", X"773", X"773", X"873", X"883", X"883", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"773", X"773", X"772", X"773", X"873", X"772", X"873", X"883", X"772", X"873", X"773", X"983", X"A94", X"983", X"983", X"A94", X"983", X"993", X"983", X"993", X"983", X"983", X"994", X"772", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"873", X"773", X"983", X"983", X"983", X"983", X"A94", X"993", X"983", X"993", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"873", X"773", X"773", X"773", X"772", X"772", X"883", X"772", X"773", X"772", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"873", X"772", X"772", X"773", X"773", X"773", X"873", X"873", X"773", X"773", X"873", X"883", X"772", X"773", X"772", X"772", X"883", X"773", X"773", X"773", X"873", X"883", X"983", X"983"),
    (X"773", X"772", X"773", X"873", X"772", X"773", X"772", X"873", X"773", X"873", X"873", X"772", X"773", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"773", X"773", X"772", X"773", X"873", X"883", X"773", X"883", X"772", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"873", X"773", X"773", X"772", X"772", X"772", X"873", X"873", X"772", X"772", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"994", X"983", X"772", X"773", X"773", X"873", X"772", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"773", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"873", X"873", X"773", X"772", X"873", X"773", X"772", X"772", X"773", X"772", X"772", X"772", X"773", X"772", X"772", X"772", X"873", X"873", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"A94", X"983", X"A94", X"983", X"983", X"983", X"993", X"983", X"993", X"773", X"772", X"883", X"772", X"773", X"773", X"773", X"883", X"773", X"773", X"772", X"772", X"773", X"773", X"773", X"873", X"773", X"873", X"773", X"883", X"772", X"873", X"984", X"983", X"A94"),
    (X"773", X"773", X"873", X"773", X"772", X"773", X"772", X"773", X"772", X"773", X"873", X"773", X"873", X"983", X"983", X"983", X"983", X"983", X"994", X"983", X"883", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"873", X"873", X"773", X"873", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"873", X"873", X"773", X"773", X"883", X"772", X"773", X"773", X"873", X"773", X"773", X"873", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"773", X"773", X"773", X"772", X"773", X"773", X"772", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"772", X"883", X"773", X"773", X"883", X"772", X"773", X"773", X"773", X"773", X"873", X"873", X"773", X"873", X"772", X"772", X"873", X"773", X"773", X"773", X"883", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"A93", X"983", X"983", X"A83", X"A83", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"772", X"773", X"883", X"773", X"773", X"772", X"772", X"772", X"773", X"772", X"873", X"873", X"773", X"883", X"773", X"773"),
    (X"872", X"872", X"772", X"772", X"772", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"983", X"A93", X"983", X"983", X"983", X"A94", X"983", X"772", X"772", X"883", X"873", X"773", X"773", X"773", X"873", X"772", X"772", X"772", X"773", X"772", X"983", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"A84", X"773", X"773", X"773", X"772", X"772", X"773", X"772", X"873", X"773", X"773", X"772", X"773", X"773", X"873", X"773", X"983", X"983", X"983", X"983", X"A83", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"883", X"773", X"772", X"772", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"873", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"A94", X"983", X"A94", X"983", X"983", X"983", X"983", X"993", X"A93", X"883", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"772", X"773", X"772", X"772", X"772", X"772"),
    (X"452", X"452", X"452", X"552", X"552", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"773", X"873", X"A94", X"983", X"983", X"A94", X"983", X"772", X"773", X"773", X"773", X"773", X"773", X"772", X"873", X"772", X"773", X"773", X"873", X"773", X"883", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"983", X"994", X"983", X"773", X"873", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"883", X"873", X"873", X"773", X"773", X"772", X"983", X"983", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"883", X"773", X"773", X"773", X"772", X"873", X"773", X"772", X"773", X"773", X"772", X"873", X"873", X"873", X"772", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"873", X"873", X"773", X"873", X"772", X"773", X"772", X"772", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"873", X"773", X"773", X"773", X"773", X"772", X"773", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"A94", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"772", X"773", X"873", X"773", X"772", X"773", X"772", X"773"),
    (X"452", X"452", X"552", X"552", X"452", X"772", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"983", X"A93", X"983", X"983", X"983", X"772", X"883", X"883", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"883", X"772", X"773", X"773", X"773", X"A94", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"773", X"873", X"883", X"883", X"772", X"773", X"772", X"772", X"772", X"772", X"773", X"773", X"772", X"873", X"773", X"983", X"994", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"772", X"883", X"883", X"873", X"873", X"772", X"773", X"773", X"772", X"773", X"773", X"772", X"883", X"873", X"773", X"983", X"993", X"A94", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"883", X"772", X"873", X"873", X"873", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"873", X"873", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"994", X"983", X"A94", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"A94", X"983", X"772", X"873", X"773", X"773", X"873", X"873", X"772", X"773", X"773", X"773"),
    (X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"772", X"773", X"773", X"773", X"773", X"883", X"883", X"773", X"773", X"772", X"883", X"772", X"773", X"773", X"873", X"983", X"983", X"983", X"983", X"A93", X"983", X"983", X"983", X"983", X"983", X"772", X"772", X"773", X"773", X"773", X"772", X"773", X"873", X"873", X"772", X"773", X"772", X"873", X"883", X"873", X"873", X"773", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"873", X"773", X"773", X"772", X"773", X"773", X"773", X"772", X"873", X"773", X"773", X"873", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"773", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"773", X"772", X"772", X"873", X"773", X"773", X"773", X"772", X"772", X"773", X"773", X"772", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"873", X"773", X"772", X"773"),
    (X"562", X"562", X"562", X"562", X"662", X"562", X"552", X"563", X"552", X"562", X"553", X"452", X"452", X"452", X"452", X"552", X"452", X"552", X"552", X"562", X"452", X"663", X"552", X"452", X"552", X"773", X"873", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"883", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"993", X"A94", X"983", X"983", X"993", X"773", X"773", X"772", X"772", X"773", X"873", X"773", X"773", X"773", X"873", X"873", X"873", X"773", X"772", X"772", X"772", X"873", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"772", X"773", X"772", X"873", X"772", X"772", X"883", X"883", X"772", X"883", X"873", X"773", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"773", X"773", X"773", X"883", X"773", X"773", X"772", X"772", X"773", X"772", X"873", X"772", X"773", X"772", X"773", X"772", X"773", X"773", X"773", X"762", X"773", X"883", X"873", X"773", X"873", X"772", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"A94", X"983", X"A94"),
    (X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"663", X"562", X"562", X"452", X"452", X"552", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"563", X"552", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"773", X"772", X"883", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"873", X"773", X"773", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"773", X"873", X"772", X"873", X"772", X"873", X"772", X"772", X"772", X"773", X"873", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"773", X"873", X"883", X"772", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"883", X"772", X"772", X"873", X"773", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"562", X"562", X"662", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"552", X"562", X"552", X"452", X"452", X"452", X"563", X"553", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"873", X"773", X"773", X"773", X"773", X"983", X"994", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"773", X"773", X"883", X"773", X"772", X"873", X"773", X"883", X"773", X"773", X"772", X"773", X"773", X"873", X"773", X"773", X"883", X"873", X"773", X"773", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"873", X"873", X"772", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"772", X"772", X"773", X"873", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"994", X"A83", X"A83", X"983", X"983", X"A94", X"773", X"772", X"772", X"873", X"773", X"883", X"773", X"873", X"773", X"773", X"772", X"773", X"773", X"873", X"772", X"773", X"772", X"773", X"772", X"773", X"773", X"772", X"873", X"772", X"772", X"773", X"773", X"772", X"773", X"873", X"993", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"662", X"562", X"452", X"452", X"452", X"552", X"452", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"773", X"873", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"773", X"773", X"772", X"772", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"873", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"773", X"773", X"773", X"773", X"773", X"772", X"883", X"873", X"772", X"772", X"873", X"773", X"773", X"773", X"772", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"883", X"772", X"772", X"883", X"772", X"773", X"773", X"773", X"883", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"A94"),
    (X"452", X"452", X"452", X"552", X"552", X"552", X"552", X"452", X"452", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"983", X"983", X"983", X"A94", X"983", X"983", X"993", X"983", X"983", X"983", X"873", X"773", X"773", X"773", X"883", X"772", X"772", X"873", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"773", X"773", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"A94", X"983", X"983", X"983", X"A93", X"983", X"983", X"983", X"772", X"773", X"772", X"772", X"772", X"772", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"773", X"873", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"772", X"772", X"773", X"773", X"772", X"873", X"773", X"772", X"773", X"873", X"773", X"772", X"772", X"773", X"873", X"773", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"772", X"883", X"773", X"873"),
    (X"452", X"452", X"552", X"452", X"452", X"552", X"452", X"452", X"563", X"452", X"552", X"562", X"662", X"562", X"562", X"562", X"662", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"883", X"772", X"773", X"772", X"772", X"773", X"772", X"773", X"772", X"773", X"773", X"883", X"873", X"773", X"773", X"773", X"772", X"773", X"772", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"A93", X"772", X"873", X"772", X"773", X"773", X"773", X"883", X"773", X"772", X"773", X"772", X"772", X"772", X"873", X"883", X"773", X"772", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"883", X"773", X"772", X"772", X"772", X"772", X"773", X"873", X"873", X"873", X"873", X"773", X"773", X"773", X"772", X"772", X"883", X"773", X"773", X"772", X"772", X"772", X"773", X"873", X"773", X"873", X"873", X"773", X"773", X"773", X"773"),
    (X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"452", X"562", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"552", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"552", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"552", X"562", X"552", X"452", X"452", X"552", X"451", X"452", X"773", X"773", X"773", X"773", X"883", X"873", X"773", X"772", X"773", X"773", X"873", X"773", X"772", X"772", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"772", X"883", X"873", X"773", X"983", X"A94", X"983", X"983", X"983", X"993", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"A94", X"773", X"873", X"773", X"772", X"773", X"773", X"772", X"773", X"772", X"873", X"873", X"773", X"873", X"772", X"873", X"873", X"773", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"773", X"773", X"773", X"773", X"773", X"883", X"773", X"773", X"773", X"772", X"773", X"883", X"772", X"772", X"873", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"772", X"773", X"773", X"772", X"773"),
    (X"562", X"562", X"673", X"562", X"562", X"562", X"662", X"562", X"562", X"662", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"552", X"452", X"552", X"552", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"452", X"552", X"552", X"563", X"452", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"883", X"772", X"772", X"773", X"773", X"772", X"772", X"873", X"772", X"883", X"773", X"772", X"772", X"773", X"773", X"773", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"A93", X"773", X"772", X"773", X"773", X"773", X"773", X"873", X"773", X"883", X"773", X"772", X"772", X"883", X"773", X"773", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"772", X"883", X"773", X"773", X"773", X"773", X"883", X"772", X"883", X"773", X"773", X"773", X"873", X"773", X"773", X"772", X"773", X"773", X"773", X"773"),
    (X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"552", X"452", X"452", X"552", X"452", X"552", X"452", X"452", X"452", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"552", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"563", X"452", X"552", X"452", X"452", X"452", X"552", X"552", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"552", X"452", X"773", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"873", X"773", X"773", X"773", X"772", X"772", X"773", X"883", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"773", X"873", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"772", X"772", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"772", X"773", X"773", X"873", X"773", X"883", X"772", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"873", X"773", X"773"),
    (X"562", X"562", X"562", X"662", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"663", X"562", X"562", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"563", X"452", X"452", X"452", X"452", X"552", X"773", X"773", X"883", X"772", X"772", X"873", X"773", X"773", X"883", X"772", X"772", X"772", X"773", X"883", X"773", X"773", X"773", X"773", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"873", X"773", X"773", X"873", X"883", X"773", X"772", X"773", X"772", X"772", X"772", X"772", X"873", X"772", X"773", X"883", X"883", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"772", X"773", X"773", X"772", X"772", X"773", X"773", X"772", X"772", X"773", X"773", X"772", X"773", X"773", X"772", X"772", X"772", X"772", X"773", X"773", X"773", X"773"),
    (X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"662", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"662", X"452", X"452", X"452", X"452", X"552", X"452", X"552", X"452", X"452", X"452", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"773", X"873", X"773", X"772", X"773", X"773", X"773", X"772", X"773", X"873", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"773", X"773", X"773", X"883", X"773", X"772", X"773", X"773", X"773", X"883", X"773", X"773", X"773", X"772", X"772", X"772", X"772", X"983", X"983", X"A94", X"983", X"A94", X"983", X"A94", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"773", X"773", X"772", X"873", X"772", X"773", X"773", X"773", X"873", X"773", X"873", X"883", X"772", X"772", X"772"),
    (X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"662", X"562", X"562", X"562", X"662", X"562", X"562", X"663", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"673", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"663", X"452", X"552", X"452", X"553", X"552", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"552", X"452", X"873", X"872", X"873", X"872", X"772", X"772", X"772", X"872", X"772", X"772", X"A83", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"994", X"983", X"983", X"A94", X"A94", X"773", X"773", X"773", X"873", X"773", X"773", X"773", X"773", X"773", X"883", X"772", X"773", X"773", X"883", X"773", X"773", X"873", X"983", X"983", X"983", X"983", X"A93", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"873", X"773", X"773", X"772", X"873", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"773", X"873", X"773"),
    (X"452", X"452", X"563", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"663", X"562", X"562", X"662", X"552", X"452", X"452", X"452", X"452", X"452", X"552", X"553", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"452", X"452", X"563", X"553", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"663", X"452", X"452", X"452", X"452", X"452", X"773", X"773", X"873", X"773", X"772", X"983", X"983", X"983", X"983", X"983", X"993", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"873", X"883", X"773", X"773", X"772", X"873", X"772", X"773", X"773", X"773", X"773", X"873", X"873", X"773", X"772", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"773", X"773", X"773", X"772", X"772", X"773", X"773", X"773", X"873", X"772", X"772", X"873"),
    (X"452", X"452", X"452", X"552", X"452", X"552", X"452", X"452", X"552", X"452", X"562", X"662", X"662", X"563", X"562", X"662", X"662", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"452", X"452", X"562", X"552", X"452", X"452", X"562", X"663", X"562", X"562", X"662", X"662", X"662", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"563", X"552", X"552", X"552", X"452", X"883", X"873", X"984", X"883", X"884", X"AA5", X"A94", X"BA5", X"AA5", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"883", X"883", X"873", X"773", X"773", X"773", X"773", X"772", X"772", X"873", X"773", X"772", X"773", X"773", X"772", X"873", X"773", X"A94", X"A94", X"993", X"A94", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"983", X"983", X"983", X"983", X"983", X"983", X"772", X"773", X"772", X"773", X"773", X"873", X"773", X"773", X"773", X"873", X"773", X"773"),
    (X"452", X"452", X"553", X"452", X"452", X"452", X"552", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"552", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"552", X"452", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"A94", X"983", X"983", X"983", X"A94", X"983", X"983", X"993", X"983", X"983", X"983", X"773", X"773", X"772", X"773", X"772", X"873", X"773", X"773", X"773", X"773", X"772", X"772", X"772", X"772", X"772", X"773", X"773", X"873", X"773", X"772", X"983", X"993", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"A83", X"873", X"773", X"772", X"773", X"773", X"772", X"773"),
    (X"673", X"562", X"552", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"452", X"452", X"452", X"552", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"562", X"552", X"552", X"562", X"552", X"552", X"552", X"552", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"562", X"562", X"673", X"663", X"562", X"663", X"552", X"562", X"552", X"562", X"552", X"452", X"552", X"552", X"562", X"552", X"563", X"452", X"552", X"552", X"662", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"563", X"562", X"562", X"562", X"663", X"552", X"552", X"562", X"452", X"452", X"452", X"452", X"452", X"663", X"452", X"452", X"452", X"452", X"563", X"452", X"563", X"552", X"552", X"552", X"552", X"562", X"563", X"562", X"563", X"562", X"983", X"983", X"A94", X"983", X"A84", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"993", X"983", X"773", X"873", X"773", X"773", X"772", X"773", X"773", X"873", X"773", X"772", X"773", X"873", X"773", X"772", X"772", X"873", X"873", X"873", X"883", X"772", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"883", X"983", X"983"),
    (X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"552", X"563", X"452", X"452", X"452", X"452", X"552", X"562", X"562", X"562", X"562", X"562", X"663", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"452", X"452", X"552", X"452", X"552", X"563", X"552", X"452", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"452", X"452", X"562", X"452", X"552", X"452", X"452", X"563", X"452", X"452", X"452", X"552", X"563", X"452", X"552", X"452", X"552", X"452", X"452", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"773", X"773", X"772", X"772", X"873", X"773", X"873", X"873", X"873", X"772", X"773", X"773", X"773", X"773", X"772", X"873", X"772", X"773", X"873", X"772", X"983", X"983", X"A94", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"994", X"983", X"983", X"983", X"983", X"983", X"983", X"994", X"983"),
    (X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"662", X"562", X"563", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"563", X"452", X"452", X"552", X"452", X"452", X"452", X"552", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"552", X"452", X"452", X"452", X"552", X"562", X"562", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"662", X"562", X"663", X"562", X"552", X"562", X"562", X"452", X"563", X"562", X"452", X"552", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"452", X"452", X"442", X"452", X"452", X"452", X"452", X"342", X"442", X"442", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"A93", X"772", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"773", X"772", X"772", X"773", X"773", X"773", X"773", X"772", X"773", X"772", X"772", X"772", X"A94", X"993", X"983", X"983", X"A94", X"983", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983"),
    (X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"552", X"552", X"563", X"452", X"452", X"452", X"452", X"552", X"563", X"452", X"562", X"662", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"662", X"662", X"562", X"562", X"673", X"663", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"663", X"562", X"562", X"562", X"562", X"553", X"452", X"452", X"452", X"452", X"562", X"562", X"562", X"562", X"562", X"673", X"562", X"562", X"562", X"562", X"552", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"562", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"452", X"563", X"452", X"452", X"663", X"452", X"452", X"452", X"552", X"552", X"452", X"452", X"452", X"983", X"983", X"983", X"A94", X"983", X"983", X"983", X"A93", X"773", X"773", X"772", X"772", X"772", X"873", X"773", X"773", X"873", X"773", X"883", X"773", X"773", X"772", X"873", X"773", X"772", X"772", X"773", X"773", X"772", X"883", X"983", X"983", X"994", X"983", X"A94", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983", X"983")
);
